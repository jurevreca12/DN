module GP_counter // General Purpose counter        
    #(parameter PRESCALER_WIDTH = 14,
      parameter LIMIT = 10000)
    (
        input logic clock,
        input logic reset,
        input start,
        output logic sample_tick
    );

    logic [PRESCALER_WIDTH-1:0] count;

    always_ff @( posedge clock) begin 
        if (reset) begin
            count <= 0;
            sample_tick <= 0;
        end
        else begin
            if (start) begin
                count <= count + 1;
                if (count == LIMIT-1) begin
                    count <= 0;
                    sample_tick <= 1;
                end
                else begin
                    sample_tick <= 0;
                end
            end 
        end
    end  
endmodule



// Components for 7-segment display

module anode_assert (
    input logic clock,
    input logic reset,
    input logic clock_enable,
    input logic enable_7seg,
    output logic [7:0] anode_select
);

    // counter that counts from 0 to 7
    logic [2:0] count;

    always_ff @(posedge clock) begin
        if (reset) begin
            count <= 0;
        end
        else begin
            if (clock_enable) begin
                count <= count + 1;
            end
        end
    end

    // assert anode_select
    assign anode_select = enable_7seg ? ~(1 << count) : ~0  ;
    
endmodule


module value_to_digit(
    input logic [31:0] value,
    input logic [7:0] anode_select,
    output logic [3:0] digit
);

    always_comb begin : value_to_digit
        case (~anode_select)
            8'H01: digit = value[3:0];
            8'H02: digit = value[7:4];
            8'H04: digit = value[11:8];
            8'H08: digit = value[15:12];
            8'H10: digit = value[19:16];
            8'H20: digit = value[23:20];
            8'H40: digit = value[27:24];
            8'H80: digit = value[31:28];
            default: digit = 4'b1111;
        endcase
    end

endmodule

// purely comb module 

module digit_to_segments (
    input logic [3:0] digit,
    output logic [6:0] segs
);
    
    always_comb begin : segDecoder
        case (digit)
            4'b0000: segs = 7'b1000000; // 0
            4'b0001: segs = 7'b1111001; // 1
            4'b0010: segs = 7'b0100100; // 2
            4'b0011: segs = 7'b0110000; // 3
            4'b0100: segs = 7'b0011001; // 4
            4'b0101: segs = 7'b0010010; // 5
            4'b0110: segs = 7'b0000010; // 6
            4'b0111: segs = 7'b1111000; // 7
            4'b1000: segs = 7'b0000000; // 8
            4'b1001: segs = 7'b0010000; // 9
            4'b1010: segs = 7'b0001000; // A
            4'b1011: segs = 7'b0000011; // b
            4'b1100: segs = 7'b1000110; // C
            4'b1101: segs = 7'b0100001; // d
            4'b1110: segs = 7'b0000110; // E
            4'b1111: segs = 7'b0001110; // F
            default: segs = 7'b1111111; // off
        endcase
    end

endmodule




module SevSegDisplay (
    input logic clock,
    input logic reset,
    input logic enable_7seg,
    input logic [3:0] digit1,
    input logic [3:0] digit2,
    input logic [3:0] digit3,
    input logic [3:0] digit4,
    input logic [3:0] digit5,
    input logic [3:0] digit6,
    input logic [3:0] digit7,
    input logic [3:0] digit8,
    output logic [7:0] anode_select,
    output logic [6:0] segs
);

    // prescaler for anode
    localparam PRESCALER_ANODE_WIDTH = 16;
    localparam PRESCALER_ANODE_LIMIT = 40000; // achieve   delay
    logic anode_clock_enable;


    // define the prescaler module for anode as GP_counter
    GP_counter #(
        .PRESCALER_WIDTH(PRESCALER_ANODE_WIDTH),
        .LIMIT(PRESCALER_ANODE_LIMIT)
    ) anode_prescaler (
        .clock(clock),
        .reset(reset),
        .start(enable_7seg),
        .sample_tick(anode_clock_enable)
    );

    // define the anode_assert module
    anode_assert anode_assert_inst (
        .clock(clock),
        .reset(reset),
        .clock_enable(anode_clock_enable),
        .enable_7seg(enable_7seg),
        .anode_select(anode_select)
    );

    // define the value_to_digit module
    logic [31:0] digit_all;
    assign digit_all = {digit8, digit7, digit6, digit5, digit4, digit3, digit2, digit1};
    logic [3:0] digit_select;

    value_to_digit value_to_digit_inst (
        .value(digit_all),
        .anode_select(anode_select),
        .digit(digit_select)
    );

    digit_to_segments digit_to_segments_inst (
        .digit(digit_select),
        .segs(segs)
    );
    
    
endmodule


`define CONFIG_REG 7'h00
`define DIGITS_REG 7'h04

module APB_7seg_display #(
    // Configurable Parameters
    parameter DW = 32 ,  // Data width
    parameter AW = 32  ,  // Address width
    // Derived Parameters
    localparam CW = 1 + DW + AW ,  // Command width  {pWRITE, pWDATA, pADDR}  
    localparam RW =  DW              // Response width { pRDATA}
)(
    input logic pCLK,
    input logic pRESETn,

    // APB signals
    input  logic [AW-1:0]  pADDR,
    input  logic           pSEL, // for each peripheral
    input  logic           pENABLE,
    input  logic           pWRITE,
    input  logic [DW-1:0]  pWDATA,
    output logic [DW-1:0]  pRDATA,
    output logic           pREADY,
    output logic           pSLVERR,

    // to fpga pins
    output logic [7:0] anode_select,
    output logic [6:0] segs
);
    // instantiate the SevSegDisplay
    logic [31:0] display_data;
    logic write_display, read_display;
    logic enable_7seg;
    logic write_config, read_config;

    SevSegDisplay SevSegDisplay_inst (
        .clock(pCLK),
        .reset(!pRESETn),
        .enable_7seg(enable_7seg), 
        .digit1(display_data[3:0]),
        .digit2(display_data[7:4]),
        .digit3(display_data[11:8]),
        .digit4(display_data[15:12]),
        .digit5(display_data[19:16]),
        .digit6(display_data[23:20]),
        .digit7(display_data[27:24]),
        .digit8(display_data[31:28]),
        .anode_select(anode_select),
        .segs(segs)
    );
    
    always_ff @(posedge pCLK) begin 
        if (!pRESETn)
            display_data <= '0;
        else if (write_display)
            display_data <= pWDATA;
    end 
    
    always_ff @(posedge pCLK) begin
        if (!pRESETn)
            enable_7seg <= 1'b0;
        else if (write_config)
            enable_7seg <= pWDATA[0]; // First bit is the enable signal
    end
    
    assign write_config  = pSEL & pWRITE & pREADY & pENABLE & pADDR[6:0] == `CONFIG_REG;
    assign write_display = pSEL & pWRITE & pREADY & pENABLE & pADDR[6:0] == `DIGITS_REG;
    assign read_config   = pSEL & !pWRITE & pREADY & pENABLE & pADDR[6:0] == `CONFIG_REG;
    assign read_display  = pSEL & !pWRITE & pREADY & pENABLE & pADDR[6:0] == `DIGITS_REG;
    
    always_comb begin
        if (read_config)
            pRDATA = {31'b0, enable_7seg};
        else if (read_display)
            pRDATA = display_data;
        else
            pRDATA = '0;
    end
    
    assign pREADY = 1'b1;
    
    logic error;
    assign error = pSEL & pREADY & pENABLE & (pADDR != `CONFIG_REG || pADDR != `DIGITS_REG);

    always_ff @(posedge pCLK) begin
        if (!pRESETn) 
            pSLVERR <= 1'b0;
        else 
            pSLVERR <= error;
    end


endmodule
